---- non-zero words: 1181
---- FILLING with 867 ----
--
-- Inferred program rom test for PicoBlaze
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity monitor is

  port (
    address     : in  std_logic_vector(11 downto 0);
    instruction : out std_logic_vector(17 downto 0);
    addr_2      : in  std_logic_vector(11 downto 0);
    wen         : in  std_logic;                    
    di          : in  std_logic_vector(17 downto 0);
    do          : out std_logic_vector(17 downto 0);
    msize       : out std_logic_vector(11 downto 0);
    clk         : in  std_logic);

end entity monitor;


architecture syn of monitor is
  -- N.B. (0 to nn) order needed otherwise data is backwards!
  type ram_type is array (0 to 2047 ) of std_logic_vector(19 downto 0);
  signal RAM : ram_type := (
    X"22020",
    X"2249C",
    X"22029",
    X"2220E",
    X"22209",
    X"22263",
    X"22249",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"0108B",
    X"2D001",
    X"01002",
    X"2D002",
    X"01A00",
    X"01C00",
    X"20288",
    X"20206",
    X"201B3",
    X"0153E",
    X"20209",
    X"01801",
    X"2020E",
    X"1D508",
    X"32045",
    X"1D50D",
    X"3204A",
    X"1D510",
    X"3203D",
    X"1D50E",
    X"32044",
    X"1D520",
    X"3A02C",
    X"1D81F",
    X"3202C",
    X"20209",
    X"2E580",
    X"11801",
    X"2202C",
    X"01880",
    X"01900",
    X"01720",
    X"2029D",
    X"01801",
    X"20282",
    X"2202C",
    X"2203D",
    X"1D801",
    X"3202C",
    X"19801",
    X"20209",
    X"2202C",
    X"2025B",
    X"01000",
    X"2E080",
    X"2F800",
    X"01980",
    X"01800",
    X"01720",
    X"2029D",
    X"01801",
    X"01A21",
    X"01B28",
    X"01C0F",
    X"20288",
    X"01A21",
    X"01900",
    X"0A080",
    X"1D000",
    X"3206A",
    X"1D020",
    X"36060",
    X"11801",
    X"22059",
    X"11901",
    X"2E8A0",
    X"11A01",
    X"00C80",
    X"0A080",
    X"11801",
    X"1D000",
    X"3206A",
    X"1D020",
    X"36064",
    X"00D80",
    X"18DC0",
    X"19D01",
    X"2EDB0",
    X"11B01",
    X"1D000",
    X"32073",
    X"1D906",
    X"36059",
    X"2F920",
    X"0B920",
    X"01A21",
    X"01B30",
    X"1D900",
    X"320A4",
    X"0A8A0",
    X"06000",
    X"06110",
    X"06220",
    X"06330",
    X"0A580",
    X"11801",
    X"1D520",
    X"32099",
    X"1D500",
    X"32099",
    X"2021A",
    X"3A087",
    X"2207E",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"14006",
    X"14100",
    X"14200",
    X"14300",
    X"04050",
    X"2207E",
    X"2E0B0",
    X"11B01",
    X"2E1B0",
    X"11B01",
    X"2E2B0",
    X"11B01",
    X"2E3B0",
    X"11B01",
    X"11A01",
    X"19901",
    X"22077",
    X"0B501",
    X"0355F",
    X"0B020",
    X"1D550",
    X"32186",
    X"1D553",
    X"3217A",
    X"1D545",
    X"3216D",
    X"1D542",
    X"32128",
    X"1D54A",
    X"32125",
    X"1D549",
    X"32108",
    X"1D54F",
    X"32117",
    X"1D552",
    X"320EE",
    X"1D557",
    X"320E7",
    X"1D554",
    X"320E3",
    X"1D548",
    X"320E1",
    X"1D543",
    X"320CA",
    X"1D556",
    X"320C5",
    X"01B01",
    X"01ACC",
    X"20249",
    X"22029",
    X"0B634",
    X"0B735",
    X"2D702",
    X"2D601",
    X"22029",
    X"01A30",
    X"01B00",
    X"2FA30",
    X"2FB31",
    X"2FB32",
    X"2FB33",
    X"01830",
    X"20103",
    X"01834",
    X"20106",
    X"01B01",
    X"2FB33",
    X"01830",
    X"20103",
    X"01838",
    X"20106",
    X"01B10",
    X"2FB33",
    X"01830",
    X"20103",
    X"01838",
    X"20106",
    X"22029",
    X"201B9",
    X"22029",
    X"0B834",
    X"0B738",
    X"2028E",
    X"2217A",
    X"1D003",
    X"360C1",
    X"01834",
    X"20103",
    X"01838",
    X"20106",
    X"22029",
    X"01A01",
    X"1D003",
    X"360F2",
    X"0BA38",
    X"01834",
    X"01704",
    X"20274",
    X"2025F",
    X"01834",
    X"20103",
    X"09007",
    X"0180C",
    X"01704",
    X"2027B",
    X"2025B",
    X"19A01",
    X"32029",
    X"01834",
    X"01704",
    X"2028E",
    X"220F2",
    X"01908",
    X"01704",
    X"22296",
    X"0190C",
    X"22104",
    X"0B734",
    X"01801",
    X"1D003",
    X"3610D",
    X"0B838",
    X"00470",
    X"20263",
    X"2025F",
    X"08470",
    X"20263",
    X"2025B",
    X"11701",
    X"19801",
    X"3610D",
    X"22029",
    X"1D003",
    X"360C1",
    X"01A38",
    X"0B82A",
    X"0B634",
    X"0A7A0",
    X"2C760",
    X"11A01",
    X"11601",
    X"19801",
    X"32029",
    X"19801",
    X"3611C",
    X"22029",
    X"0B634",
    X"0B735",
    X"26760",
    X"2020E",
    X"00650",
    X"1D62B",
    X"32139",
    X"1D63D",
    X"3213E",
    X"1D624",
    X"36128",
    X"20148",
    X"360C1",
    X"00470",
    X"20263",
    X"00460",
    X"20137",
    X"22029",
    X"20263",
    X"2225B",
    X"20148",
    X"360C1",
    X"00A60",
    X"00B70",
    X"22128",
    X"20148",
    X"360C1",
    X"2DA03",
    X"2DB04",
    X"2D605",
    X"2D706",
    X"2D807",
    X"11A01",
    X"13B00",
    X"22128",
    X"20164",
    X"35000",
    X"00840",
    X"1480E",
    X"1480E",
    X"1480E",
    X"1480E",
    X"00740",
    X"14706",
    X"14706",
    X"14706",
    X"14706",
    X"20164",
    X"35000",
    X"00540",
    X"1450E",
    X"1450E",
    X"04750",
    X"1440C",
    X"1440C",
    X"01600",
    X"04640",
    X"036C0",
    X"20164",
    X"35000",
    X"04640",
    X"06000",
    X"25000",
    X"2020E",
    X"19520",
    X"39000",
    X"1D540",
    X"3D000",
    X"0353F",
    X"00450",
    X"06000",
    X"25000",
    X"1D003",
    X"360C1",
    X"0B634",
    X"0B735",
    X"2D603",
    X"2D704",
    X"0B638",
    X"2D605",
    X"0B639",
    X"2D606",
    X"0B63A",
    X"2D607",
    X"22029",
    X"01600",
    X"0187F",
    X"1D002",
    X"3A183",
    X"0B634",
    X"1D003",
    X"3A183",
    X"0B838",
    X"19801",
    X"201A5",
    X"2025B",
    X"22029",
    X"01600",
    X"01700",
    X"01810",
    X"1D002",
    X"3A190",
    X"0B634",
    X"0B735",
    X"1D003",
    X"3A190",
    X"0B838",
    X"20192",
    X"22029",
    X"2D603",
    X"2D704",
    X"00470",
    X"20263",
    X"00460",
    X"20263",
    X"2025F",
    X"09405",
    X"20263",
    X"09404",
    X"20263",
    X"09403",
    X"20263",
    X"2025B",
    X"11601",
    X"13700",
    X"19801",
    X"3A029",
    X"22192",
    X"00460",
    X"20263",
    X"2025F",
    X"2025F",
    X"0A460",
    X"20263",
    X"2025F",
    X"11601",
    X"19801",
    X"39000",
    X"0D60F",
    X"361A9",
    X"2025B",
    X"221A5",
    X"01B01",
    X"01ABD",
    X"20249",
    X"14580",
    X"20209",
    X"25000",
    X"01B02",
    X"01AA4",
    X"20250",
    X"25000",
    X"2154D",
    X"2156F",
    X"2156E",
    X"21569",
    X"21574",
    X"2156F",
    X"21572",
    X"21520",
    X"21556",
    X"21532",
    X"2152E",
    X"21531",
    X"2150D",
    X"2150A",
    X"21500",
    X"21545",
    X"21572",
    X"21572",
    X"2156F",
    X"21572",
    X"2150D",
    X"2150A",
    X"21500",
    X"21553",
    X"21520",
    X"2155B",
    X"21528",
    X"21573",
    X"21574",
    X"21561",
    X"21572",
    X"21574",
    X"21529",
    X"21520",
    X"2155B",
    X"21528",
    X"21563",
    X"2156F",
    X"21575",
    X"2156E",
    X"21574",
    X"21529",
    X"2155D",
    X"2155D",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21564",
    X"21575",
    X"2156D",
    X"21570",
    X"21520",
    X"21573",
    X"21563",
    X"21572",
    X"21561",
    X"21574",
    X"21563",
    X"21568",
    X"21570",
    X"21561",
    X"21564",
    X"21520",
    X"2156D",
    X"21565",
    X"2156D",
    X"2156F",
    X"21572",
    X"21579",
    X"21524",
    X"21500",
    X"2B031",
    X"2B001",
    X"25000",
    X"09000",
    X"0D004",
    X"36209",
    X"2D580",
    X"25000",
    X"20211",
    X"35000",
    X"2220E",
    X"011A7",
    X"09000",
    X"0D008",
    X"36218",
    X"19101",
    X"31000",
    X"22212",
    X"09501",
    X"25000",
    X"19530",
    X"3A228",
    X"1D50A",
    X"3A22B",
    X"19511",
    X"3A228",
    X"1150A",
    X"1D510",
    X"3A22B",
    X"1952A",
    X"3A228",
    X"1150A",
    X"1D510",
    X"3A22B",
    X"01500",
    X"1450E",
    X"25000",
    X"25000",
    X"2020E",
    X"20209",
    X"2021A",
    X"39000",
    X"01507",
    X"20209",
    X"2222C",
    X"00510",
    X"2021A",
    X"3D000",
    X"00450",
    X"14406",
    X"14406",
    X"14406",
    X"14406",
    X"00500",
    X"2021A",
    X"3D000",
    X"04450",
    X"25000",
    X"2022C",
    X"00450",
    X"14406",
    X"14406",
    X"14406",
    X"14406",
    X"2022C",
    X"04450",
    X"25000",
    X"24BA0",
    X"1D500",
    X"31000",
    X"20209",
    X"11A01",
    X"13B00",
    X"22249",
    X"24BA0",
    X"1D500",
    X"31000",
    X"1D524",
    X"36257",
    X"2025B",
    X"22258",
    X"20209",
    X"11A01",
    X"13B00",
    X"22250",
    X"0150D",
    X"20209",
    X"0150A",
    X"22209",
    X"01520",
    X"22209",
    X"11530",
    X"22209",
    X"00540",
    X"1450E",
    X"1450E",
    X"1450E",
    X"1450E",
    X"2026F",
    X"20209",
    X"00540",
    X"0350F",
    X"2026F",
    X"20209",
    X"25000",
    X"1950A",
    X"3A272",
    X"11507",
    X"1153A",
    X"25000",
    X"10870",
    X"19801",
    X"0A480",
    X"20263",
    X"19701",
    X"31000",
    X"22275",
    X"10870",
    X"19801",
    X"08480",
    X"20263",
    X"19701",
    X"31000",
    X"2227C",
    X"0A580",
    X"04550",
    X"31000",
    X"20209",
    X"11801",
    X"22282",
    X"01900",
    X"2E9A0",
    X"11A01",
    X"19C01",
    X"36288",
    X"25000",
    X"0A080",
    X"11001",
    X"2E080",
    X"3D000",
    X"11801",
    X"19701",
    X"3628E",
    X"25000",
    X"0A080",
    X"2C090",
    X"11801",
    X"11901",
    X"19701",
    X"36296",
    X"25000",
    X"0A080",
    X"2E090",
    X"11801",
    X"11901",
    X"19701",
    X"3629D",
    X"25000",
    X"21553",
    X"21520",
    X"2155B",
    X"21528",
    X"21573",
    X"21574",
    X"21561",
    X"21572",
    X"21574",
    X"21529",
    X"21520",
    X"2155B",
    X"21528",
    X"21563",
    X"2156F",
    X"21575",
    X"2156E",
    X"21574",
    X"21529",
    X"2155D",
    X"2155D",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21564",
    X"21575",
    X"2156D",
    X"21570",
    X"21520",
    X"21573",
    X"21563",
    X"21572",
    X"21561",
    X"21574",
    X"21563",
    X"21568",
    X"21570",
    X"21561",
    X"21564",
    X"21520",
    X"2156D",
    X"21565",
    X"2156D",
    X"2156F",
    X"21572",
    X"21579",
    X"21524",
    X"21570",
    X"21520",
    X"2155B",
    X"21528",
    X"21573",
    X"21574",
    X"21561",
    X"21572",
    X"21574",
    X"21529",
    X"21520",
    X"2155B",
    X"21528",
    X"21563",
    X"2156F",
    X"21575",
    X"2156E",
    X"21574",
    X"21529",
    X"2155D",
    X"2155D",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21564",
    X"21575",
    X"2156D",
    X"21570",
    X"21520",
    X"21570",
    X"21572",
    X"2156F",
    X"21567",
    X"21572",
    X"21561",
    X"2156D",
    X"21520",
    X"2156D",
    X"21565",
    X"2156D",
    X"2156F",
    X"21572",
    X"21579",
    X"21524",
    X"21565",
    X"21520",
    X"21528",
    X"21561",
    X"21564",
    X"21564",
    X"21572",
    X"21529",
    X"21520",
    X"21528",
    X"21564",
    X"21561",
    X"21574",
    X"21561",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21565",
    X"21564",
    X"21569",
    X"21574",
    X"21520",
    X"21570",
    X"21572",
    X"2156F",
    X"21567",
    X"21572",
    X"21561",
    X"2156D",
    X"21520",
    X"2156D",
    X"21565",
    X"2156D",
    X"2156F",
    X"21572",
    X"21579",
    X"21520",
    X"21528",
    X"2156F",
    X"2156E",
    X"21565",
    X"21520",
    X"21577",
    X"2156F",
    X"21572",
    X"21564",
    X"21529",
    X"21524",
    X"21569",
    X"21520",
    X"21528",
    X"21570",
    X"2156F",
    X"21572",
    X"21574",
    X"21529",
    X"21520",
    X"2155B",
    X"21528",
    X"21563",
    X"2156F",
    X"21575",
    X"2156E",
    X"21574",
    X"21529",
    X"2155D",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21572",
    X"21565",
    X"21561",
    X"21564",
    X"21520",
    X"21549",
    X"2152F",
    X"2154F",
    X"21520",
    X"21570",
    X"2156F",
    X"21572",
    X"21574",
    X"21528",
    X"21573",
    X"21529",
    X"21524",
    X"2156F",
    X"21520",
    X"21528",
    X"21570",
    X"2156F",
    X"21572",
    X"21574",
    X"21529",
    X"21520",
    X"21528",
    X"21564",
    X"21561",
    X"21574",
    X"21561",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21577",
    X"21572",
    X"21569",
    X"21574",
    X"21565",
    X"21520",
    X"21549",
    X"2152F",
    X"2154F",
    X"21520",
    X"21570",
    X"2156F",
    X"21572",
    X"21574",
    X"21524",
    X"2156A",
    X"21520",
    X"21528",
    X"21561",
    X"21564",
    X"21564",
    X"21572",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"2156A",
    X"21575",
    X"2156D",
    X"21570",
    X"21520",
    X"21574",
    X"2156F",
    X"21520",
    X"21561",
    X"21564",
    X"21564",
    X"21572",
    X"21565",
    X"21573",
    X"21573",
    X"21524",
    X"21577",
    X"21520",
    X"21528",
    X"21561",
    X"21564",
    X"21564",
    X"21572",
    X"21529",
    X"21520",
    X"21528",
    X"21564",
    X"21561",
    X"21574",
    X"21561",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21577",
    X"21572",
    X"21569",
    X"21574",
    X"21565",
    X"21520",
    X"21574",
    X"2156F",
    X"21520",
    X"21565",
    X"2152D",
    X"21562",
    X"21575",
    X"21573",
    X"21524",
    X"21572",
    X"21520",
    X"21528",
    X"21561",
    X"21564",
    X"21564",
    X"21572",
    X"21529",
    X"21520",
    X"2155B",
    X"21528",
    X"21563",
    X"2156F",
    X"21575",
    X"2156E",
    X"21574",
    X"21529",
    X"2155D",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21572",
    X"21565",
    X"21561",
    X"21564",
    X"21520",
    X"21566",
    X"21572",
    X"2156F",
    X"2156D",
    X"21520",
    X"21565",
    X"2152D",
    X"21562",
    X"21575",
    X"21573",
    X"21524",
    X"21562",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21573",
    X"21574",
    X"21561",
    X"21572",
    X"21574",
    X"21520",
    X"21555",
    X"21555",
    X"21545",
    X"21520",
    X"21562",
    X"2156F",
    X"2156F",
    X"21574",
    X"2156C",
    X"2156F",
    X"21561",
    X"21564",
    X"21565",
    X"21572",
    X"21524",
    X"21563",
    X"21520",
    X"21528",
    X"21564",
    X"21561",
    X"21574",
    X"21561",
    X"21529",
    X"21520",
    X"21528",
    X"2156C",
    X"21565",
    X"2156E",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21577",
    X"21572",
    X"21569",
    X"21574",
    X"21565",
    X"21520",
    X"21543",
    X"21549",
    X"21554",
    X"21549",
    X"21552",
    X"2154F",
    X"21543",
    X"21520",
    X"21573",
    X"21565",
    X"21572",
    X"21569",
    X"21561",
    X"2156C",
    X"21524",
    X"21576",
    X"21520",
    X"21528",
    X"21564",
    X"21569",
    X"21576",
    X"21529",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"21520",
    X"2152D",
    X"21520",
    X"21573",
    X"21565",
    X"21574",
    X"21520",
    X"21562",
    X"21561",
    X"21575",
    X"21564",
    X"21520",
    X"21572",
    X"21561",
    X"21574",
    X"21565",
    X"21520",
    X"21564",
    X"21569",
    X"21556",
    X"21569",
    X"21573",
    X"2156F",
    X"21572",
    X"21524",
    X"21500",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000",
    X"00000"
    );
begin

  process (clk) is
  begin  -- process
    if clk'event and clk = '1' then     -- rising clock edge
      instruction <= RAM(to_integer(unsigned(address)))(17 downto 0);
      if wen = '1' then
        RAM(to_integer(unsigned(addr_2))) <= B"00" & di;
      end if;
    end if;
  end process;

  do <= RAM(to_integer(unsigned(addr_2)))(17 downto 0);

  msize <= std_logic_vector( to_unsigned( RAM'length, msize'length));

end syn;
